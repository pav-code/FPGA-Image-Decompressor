library verilog;
use verilog.vl_types.all;
entity mil1_FSM_v_unit is
end mil1_FSM_v_unit;

library verilog;
use verilog.vl_types.all;
entity mil2_FSM_v_unit is
end mil2_FSM_v_unit;
